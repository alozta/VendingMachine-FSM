library verilog;
use verilog.vl_types.all;
entity vending_machine_testbench is
end vending_machine_testbench;
